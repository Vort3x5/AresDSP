module rom_input (
    input  [11:0] addr,
    output reg signed [15:0] data_real,
    output reg signed [15:0] data_imag
);
    always @(*) begin
        case (addr)		
		12'd0   : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd1   : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd2   : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd3   : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd4   : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd5   : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd6   : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd7   : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd8   : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd9   : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd10  : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd11  : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd12  : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd13  : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd14  : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd15  : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd16  : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd17  : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd18  : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd19  : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd20  : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd21  : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd22  : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd23  : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd24  : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd25  : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd26  : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd27  : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd28  : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd29  : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd30  : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd31  : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd32  : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd33  : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd34  : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd35  : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd36  : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd37  : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd38  : begin data_real = 16'sd25088; data_imag = 16'sd0; end
		12'd39  : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd40  : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd41  : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd42  : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd43  : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd44  : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd45  : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd46  : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd47  : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd48  : begin data_real = -16'sd17664; data_imag = 16'sd0; end
		12'd49  : begin data_real = -16'sd15872; data_imag = 16'sd0; end
		12'd50  : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd51  : begin data_real = -16'sd16384; data_imag = 16'sd0; end
		12'd52  : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd53  : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd54  : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd55  : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd56  : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd57  : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd58  : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd59  : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd60  : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd61  : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd62  : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd63  : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd64  : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd65  : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd66  : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd67  : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd68  : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd69  : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd70  : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd71  : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd72  : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd73  : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd74  : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd75  : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd76  : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd77  : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd78  : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd79  : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd80  : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd81  : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd82  : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd83  : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd84  : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd85  : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd86  : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd87  : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd88  : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd89  : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd90  : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd91  : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd92  : begin data_real = 16'sd15104; data_imag = 16'sd0; end
		12'd93  : begin data_real = 16'sd16640; data_imag = 16'sd0; end
		12'd94  : begin data_real = 16'sd20480; data_imag = 16'sd0; end
		12'd95  : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd96  : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd97  : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd98  : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd99  : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd100 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd101 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd102 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd103 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd104 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd105 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd106 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd107 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd108 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd109 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd110 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd111 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd112 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd113 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd114 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd115 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd116 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd117 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd118 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd119 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd120 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd121 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd122 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd123 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd124 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd125 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd126 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd127 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd128 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd129 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd130 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd131 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd132 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd133 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd134 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd135 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd136 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd137 : begin data_real = -16'sd16640; data_imag = 16'sd0; end
		12'd138 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd139 : begin data_real = -16'sd16896; data_imag = 16'sd0; end
		12'd140 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd141 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd142 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd143 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd144 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd145 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd146 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd147 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd148 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd149 : begin data_real = 16'sd16128; data_imag = 16'sd0; end
		12'd150 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd151 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd152 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd153 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd154 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd155 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd156 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd157 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd158 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd159 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd160 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd161 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd162 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd163 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd164 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd165 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd166 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd167 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd168 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd169 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd170 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd171 : begin data_real = -16'sd17152; data_imag = 16'sd0; end
		12'd172 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd173 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd174 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd175 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd176 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd177 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd178 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd179 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd180 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd181 : begin data_real = 16'sd16128; data_imag = 16'sd0; end
		12'd182 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd183 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd184 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd185 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd186 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd187 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd188 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd189 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd190 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd191 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd192 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd193 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd194 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd195 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd196 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd197 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd198 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd199 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd200 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd201 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd202 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd203 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd204 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd205 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd206 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd207 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd208 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd209 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd210 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd211 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd212 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd213 : begin data_real = 16'sd15360; data_imag = 16'sd0; end
		12'd214 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd215 : begin data_real = 16'sd17152; data_imag = 16'sd0; end
		12'd216 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd217 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd218 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd219 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd220 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd221 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd222 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd223 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd224 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd225 : begin data_real = -16'sd16128; data_imag = 16'sd0; end
		12'd226 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd227 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd228 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd229 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd230 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd231 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd232 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd233 : begin data_real = 16'sd17152; data_imag = 16'sd0; end
		12'd234 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd235 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd236 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd237 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd238 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd239 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd240 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd241 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd242 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd243 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd244 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd245 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd246 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd247 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd248 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd249 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd250 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd251 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd252 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd253 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd254 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd255 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd256 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd257 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd258 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd259 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd260 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd261 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd262 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd263 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd264 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd265 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd266 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd267 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd268 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd269 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd270 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd271 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd272 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd273 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd274 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd275 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd276 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd277 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd278 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd279 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd280 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd281 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd282 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd283 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd284 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd285 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd286 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd287 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd288 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd289 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd290 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd291 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd292 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd293 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd294 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd295 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd296 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd297 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd298 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd299 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd300 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd301 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd302 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd303 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd304 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd305 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd306 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd307 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd308 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd309 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd310 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd311 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd312 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd313 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd314 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd315 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd316 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd317 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd318 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd319 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd320 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd321 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd322 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd323 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd324 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd325 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd326 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd327 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd328 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd329 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd330 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd331 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd332 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd333 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd334 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd335 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd336 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd337 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd338 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd339 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd340 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd341 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd342 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd343 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd344 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd345 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd346 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd347 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd348 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd349 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd350 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd351 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd352 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd353 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd354 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd355 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd356 : begin data_real = 16'sd16640; data_imag = 16'sd0; end
		12'd357 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd358 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd359 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd360 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd361 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd362 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd363 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd364 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd365 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd366 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd367 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd368 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd369 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd370 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd371 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd372 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd373 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd374 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd375 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd376 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd377 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd378 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd379 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd380 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd381 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd382 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd383 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd384 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd385 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd386 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd387 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd388 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd389 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd390 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd391 : begin data_real = 16'sd14336; data_imag = 16'sd0; end
		12'd392 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd393 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd394 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd395 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd396 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd397 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd398 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd399 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd400 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd401 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd402 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd403 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd404 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd405 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd406 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd407 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd408 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd409 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd410 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd411 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd412 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd413 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd414 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd415 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd416 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd417 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd418 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd419 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd420 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd421 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd422 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd423 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd424 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd425 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd426 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd427 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd428 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd429 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd430 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd431 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd432 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd433 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd434 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd435 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd436 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd437 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd438 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd439 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd440 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd441 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd442 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd443 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd444 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd445 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd446 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd447 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd448 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd449 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd450 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd451 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd452 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd453 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd454 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd455 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd456 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd457 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd458 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd459 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd460 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd461 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd462 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd463 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd464 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd465 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd466 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd467 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd468 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd469 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd470 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd471 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd472 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd473 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd474 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd475 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd476 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd477 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd478 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd479 : begin data_real = 16'sd15104; data_imag = 16'sd0; end
		12'd480 : begin data_real = 16'sd18432; data_imag = 16'sd0; end
		12'd481 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd482 : begin data_real = 16'sd15360; data_imag = 16'sd0; end
		12'd483 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd484 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd485 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd486 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd487 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd488 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd489 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd490 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd491 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd492 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd493 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd494 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd495 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd496 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd497 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd498 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd499 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd500 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd501 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd502 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd503 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd504 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd505 : begin data_real = -16'sd12032; data_imag = 16'sd0; end
		12'd506 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd507 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd508 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd509 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd510 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd511 : begin data_real = 16'sd15616; data_imag = 16'sd0; end
		12'd512 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd513 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd514 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd515 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd516 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd517 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd518 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd519 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd520 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd521 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd522 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd523 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd524 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd525 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd526 : begin data_real = -16'sd16896; data_imag = 16'sd0; end
		12'd527 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd528 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd529 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd530 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd531 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd532 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd533 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd534 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd535 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd536 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd537 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd538 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd539 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd540 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd541 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd542 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd543 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd544 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd545 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd546 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd547 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd548 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd549 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd550 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd551 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd552 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd553 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd554 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd555 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd556 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd557 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd558 : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd559 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd560 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd561 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd562 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd563 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd564 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd565 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd566 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd567 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd568 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd569 : begin data_real = 16'sd17920; data_imag = 16'sd0; end
		12'd570 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd571 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd572 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd573 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd574 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd575 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd576 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd577 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd578 : begin data_real = -16'sd14336; data_imag = 16'sd0; end
		12'd579 : begin data_real = -16'sd14080; data_imag = 16'sd0; end
		12'd580 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd581 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd582 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd583 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd584 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd585 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd586 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd587 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd588 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd589 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd590 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd591 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd592 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd593 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd594 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd595 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd596 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd597 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd598 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd599 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd600 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd601 : begin data_real = 16'sd16128; data_imag = 16'sd0; end
		12'd602 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd603 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd604 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd605 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd606 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd607 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd608 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd609 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd610 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd611 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd612 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd613 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd614 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd615 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd616 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd617 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd618 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd619 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd620 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd621 : begin data_real = 16'sd18176; data_imag = 16'sd0; end
		12'd622 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd623 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd624 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd625 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd626 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd627 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd628 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd629 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd630 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd631 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd632 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd633 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd634 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd635 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd636 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd637 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd638 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd639 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd640 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd641 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd642 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd643 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd644 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd645 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd646 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd647 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd648 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd649 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd650 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd651 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd652 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd653 : begin data_real = 16'sd17152; data_imag = 16'sd0; end
		12'd654 : begin data_real = 16'sd21504; data_imag = 16'sd0; end
		12'd655 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd656 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd657 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd658 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd659 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd660 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd661 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd662 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd663 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd664 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd665 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd666 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd667 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd668 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd669 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd670 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd671 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd672 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd673 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd674 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd675 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd676 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd677 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd678 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd679 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd680 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd681 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd682 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd683 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd684 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd685 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd686 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd687 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd688 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd689 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd690 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd691 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd692 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd693 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd694 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd695 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd696 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd697 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd698 : begin data_real = -16'sd18432; data_imag = 16'sd0; end
		12'd699 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd700 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd701 : begin data_real = -16'sd12032; data_imag = 16'sd0; end
		12'd702 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd703 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd704 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd705 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd706 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd707 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd708 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd709 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd710 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd711 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd712 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd713 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd714 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd715 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd716 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd717 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd718 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd719 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd720 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd721 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd722 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd723 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd724 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd725 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd726 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd727 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd728 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd729 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd730 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd731 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd732 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd733 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd734 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd735 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd736 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd737 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd738 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd739 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd740 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd741 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd742 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd743 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd744 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd745 : begin data_real = 16'sd16128; data_imag = 16'sd0; end
		12'd746 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd747 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd748 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd749 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd750 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd751 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd752 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd753 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd754 : begin data_real = -16'sd22016; data_imag = 16'sd0; end
		12'd755 : begin data_real = -16'sd15872; data_imag = 16'sd0; end
		12'd756 : begin data_real = -16'sd14336; data_imag = 16'sd0; end
		12'd757 : begin data_real = -16'sd15872; data_imag = 16'sd0; end
		12'd758 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd759 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd760 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd761 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd762 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd763 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd764 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd765 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd766 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd767 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd768 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd769 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd770 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd771 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd772 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd773 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd774 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd775 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd776 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd777 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd778 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd779 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd780 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd781 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd782 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd783 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd784 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd785 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd786 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd787 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd788 : begin data_real = -16'sd15872; data_imag = 16'sd0; end
		12'd789 : begin data_real = -16'sd22272; data_imag = 16'sd0; end
		12'd790 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd791 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd792 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd793 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd794 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd795 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd796 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd797 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd798 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd799 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd800 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd801 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd802 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd803 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd804 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd805 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd806 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd807 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd808 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd809 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd810 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd811 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd812 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd813 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd814 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd815 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd816 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd817 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd818 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd819 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd820 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd821 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd822 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd823 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd824 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd825 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd826 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd827 : begin data_real = 16'sd19200; data_imag = 16'sd0; end
		12'd828 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd829 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd830 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd831 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd832 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd833 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd834 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd835 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd836 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd837 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd838 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd839 : begin data_real = -16'sd16896; data_imag = 16'sd0; end
		12'd840 : begin data_real = -16'sd15616; data_imag = 16'sd0; end
		12'd841 : begin data_real = -16'sd17920; data_imag = 16'sd0; end
		12'd842 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd843 : begin data_real = -16'sd21248; data_imag = 16'sd0; end
		12'd844 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd845 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd846 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd847 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd848 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd849 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd850 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd851 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd852 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd853 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd854 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd855 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd856 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd857 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd858 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd859 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd860 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd861 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd862 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd863 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd864 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd865 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd866 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd867 : begin data_real = 16'sd15360; data_imag = 16'sd0; end
		12'd868 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd869 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd870 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd871 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd872 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd873 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd874 : begin data_real = -16'sd17408; data_imag = 16'sd0; end
		12'd875 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd876 : begin data_real = -16'sd18944; data_imag = 16'sd0; end
		12'd877 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd878 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd879 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd880 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd881 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd882 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd883 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd884 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd885 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd886 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd887 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd888 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd889 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd890 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd891 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd892 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd893 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd894 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd895 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd896 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd897 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd898 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd899 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd900 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd901 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd902 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd903 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd904 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd905 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd906 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd907 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd908 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd909 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd910 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd911 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd912 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd913 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd914 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd915 : begin data_real = 16'sd18688; data_imag = 16'sd0; end
		12'd916 : begin data_real = 16'sd18688; data_imag = 16'sd0; end
		12'd917 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd918 : begin data_real = 16'sd16896; data_imag = 16'sd0; end
		12'd919 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd920 : begin data_real = 16'sd18432; data_imag = 16'sd0; end
		12'd921 : begin data_real = 16'sd21504; data_imag = 16'sd0; end
		12'd922 : begin data_real = 16'sd18176; data_imag = 16'sd0; end
		12'd923 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd924 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd925 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd926 : begin data_real = -16'sd14336; data_imag = 16'sd0; end
		12'd927 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd928 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd929 : begin data_real = -16'sd24064; data_imag = 16'sd0; end
		12'd930 : begin data_real = -16'sd15872; data_imag = 16'sd0; end
		12'd931 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd932 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd933 : begin data_real = -16'sd12032; data_imag = 16'sd0; end
		12'd934 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd935 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd936 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd937 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd938 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd939 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd940 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd941 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd942 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd943 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd944 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd945 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd946 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd947 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd948 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd949 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd950 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd951 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd952 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd953 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd954 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd955 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd956 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd957 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd958 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd959 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd960 : begin data_real = -16'sd12032; data_imag = 16'sd0; end
		12'd961 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd962 : begin data_real = -16'sd18176; data_imag = 16'sd0; end
		12'd963 : begin data_real = -16'sd18176; data_imag = 16'sd0; end
		12'd964 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd965 : begin data_real = -16'sd18944; data_imag = 16'sd0; end
		12'd966 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd967 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd968 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd969 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd970 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd971 : begin data_real = 16'sd15360; data_imag = 16'sd0; end
		12'd972 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd973 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd974 : begin data_real = 16'sd16384; data_imag = 16'sd0; end
		12'd975 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd976 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd977 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd978 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd979 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd980 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd981 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd982 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd983 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd984 : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd985 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd986 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd987 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd988 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd989 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd990 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd991 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd992 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd993 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd994 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd995 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd996 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd997 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd998 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd999 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1000 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1001 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd1002 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1003 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1004 : begin data_real = 16'sd15872; data_imag = 16'sd0; end
		12'd1005 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd1006 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1007 : begin data_real = 16'sd16384; data_imag = 16'sd0; end
		12'd1008 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd1009 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1010 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1011 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1012 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1013 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1014 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd1015 : begin data_real = -16'sd18432; data_imag = 16'sd0; end
		12'd1016 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd1017 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd1018 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd1019 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd1020 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd1021 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd1022 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1023 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd1024 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd1025 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1026 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd1027 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd1028 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd1029 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1030 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd1031 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd1032 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1033 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1034 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1035 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd1036 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd1037 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1038 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1039 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1040 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd1041 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd1042 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd1043 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd1044 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd1045 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd1046 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd1047 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1048 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1049 : begin data_real = -16'sd17920; data_imag = 16'sd0; end
		12'd1050 : begin data_real = -16'sd17920; data_imag = 16'sd0; end
		12'd1051 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1052 : begin data_real = -16'sd12032; data_imag = 16'sd0; end
		12'd1053 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd1054 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1055 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1056 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd1057 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1058 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd1059 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd1060 : begin data_real = 16'sd15872; data_imag = 16'sd0; end
		12'd1061 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1062 : begin data_real = 16'sd16896; data_imag = 16'sd0; end
		12'd1063 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1064 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1065 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1066 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1067 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1068 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd1069 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1070 : begin data_real = -16'sd14080; data_imag = 16'sd0; end
		12'd1071 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd1072 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1073 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1074 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1075 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd1076 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd1077 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd1078 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1079 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd1080 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1081 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd1082 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1083 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd1084 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1085 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1086 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1087 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1088 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd1089 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1090 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1091 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1092 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd1093 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1094 : begin data_real = 16'sd17920; data_imag = 16'sd0; end
		12'd1095 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd1096 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd1097 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1098 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1099 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1100 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1101 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd1102 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd1103 : begin data_real = -16'sd20736; data_imag = 16'sd0; end
		12'd1104 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd1105 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd1106 : begin data_real = -16'sd17152; data_imag = 16'sd0; end
		12'd1107 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1108 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1109 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1110 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1111 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1112 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1113 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1114 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd1115 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1116 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd1117 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd1118 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1119 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd1120 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1121 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd1122 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1123 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1124 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1125 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd1126 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1127 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1128 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1129 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1130 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1131 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1132 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd1133 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1134 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd1135 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1136 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1137 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd1138 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd1139 : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd1140 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd1141 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1142 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd1143 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd1144 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1145 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1146 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1147 : begin data_real = 16'sd18944; data_imag = 16'sd0; end
		12'd1148 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd1149 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1150 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1151 : begin data_real = 16'sd16128; data_imag = 16'sd0; end
		12'd1152 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd1153 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1154 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1155 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd1156 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd1157 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd1158 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd1159 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1160 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd1161 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd1162 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1163 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1164 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd1165 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1166 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1167 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1168 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd1169 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1170 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd1171 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1172 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1173 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1174 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd1175 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd1176 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1177 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1178 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1179 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd1180 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1181 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1182 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd1183 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1184 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1185 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1186 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1187 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd1188 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1189 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd1190 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1191 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1192 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd1193 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd1194 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd1195 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd1196 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd1197 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1198 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1199 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1200 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1201 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1202 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1203 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd1204 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd1205 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd1206 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1207 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1208 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1209 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1210 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1211 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1212 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd1213 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1214 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1215 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1216 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd1217 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1218 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1219 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1220 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd1221 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1222 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1223 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1224 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd1225 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1226 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd1227 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd1228 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd1229 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd1230 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1231 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1232 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd1233 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1234 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1235 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1236 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd1237 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1238 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1239 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1240 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1241 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd1242 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd1243 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd1244 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1245 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd1246 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd1247 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1248 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd1249 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1250 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1251 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1252 : begin data_real = 16'sd15872; data_imag = 16'sd0; end
		12'd1253 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1254 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1255 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1256 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd1257 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1258 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd1259 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1260 : begin data_real = -16'sd16384; data_imag = 16'sd0; end
		12'd1261 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1262 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd1263 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1264 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd1265 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1266 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1267 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd1268 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd1269 : begin data_real = 16'sd15616; data_imag = 16'sd0; end
		12'd1270 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1271 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd1272 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1273 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd1274 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd1275 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1276 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1277 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1278 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd1279 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd1280 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1281 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd1282 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd1283 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd1284 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1285 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd1286 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1287 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1288 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1289 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1290 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd1291 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1292 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1293 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd1294 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd1295 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd1296 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1297 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd1298 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1299 : begin data_real = -16'sd17920; data_imag = 16'sd0; end
		12'd1300 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd1301 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1302 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1303 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd1304 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1305 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd1306 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd1307 : begin data_real = 16'sd14336; data_imag = 16'sd0; end
		12'd1308 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1309 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1310 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd1311 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd1312 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1313 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd1314 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1315 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd1316 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1317 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd1318 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd1319 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1320 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd1321 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd1322 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1323 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd1324 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd1325 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd1326 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1327 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd1328 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1329 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1330 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1331 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1332 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1333 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1334 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1335 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1336 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1337 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1338 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd1339 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1340 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1341 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1342 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1343 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1344 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1345 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1346 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1347 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1348 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd1349 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1350 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1351 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1352 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd1353 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1354 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1355 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd1356 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd1357 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd1358 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1359 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd1360 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd1361 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd1362 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1363 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1364 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1365 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1366 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1367 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1368 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1369 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1370 : begin data_real = -16'sd19200; data_imag = 16'sd0; end
		12'd1371 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1372 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1373 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1374 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1375 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1376 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1377 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd1378 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1379 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1380 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd1381 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1382 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1383 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd1384 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd1385 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1386 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1387 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1388 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd1389 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1390 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd1391 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1392 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1393 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1394 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd1395 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1396 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1397 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1398 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1399 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1400 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd1401 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1402 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1403 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd1404 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd1405 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1406 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1407 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd1408 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1409 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1410 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1411 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1412 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1413 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd1414 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1415 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1416 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1417 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1418 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1419 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd1420 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1421 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd1422 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd1423 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd1424 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1425 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1426 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd1427 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1428 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd1429 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1430 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd1431 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd1432 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1433 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd1434 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd1435 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1436 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd1437 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd1438 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1439 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd1440 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd1441 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1442 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1443 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1444 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd1445 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1446 : begin data_real = 16'sd22528; data_imag = 16'sd0; end
		12'd1447 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1448 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1449 : begin data_real = 16'sd16384; data_imag = 16'sd0; end
		12'd1450 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd1451 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1452 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd1453 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd1454 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd1455 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd1456 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1457 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd1458 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1459 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1460 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1461 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1462 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1463 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1464 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1465 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1466 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1467 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1468 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1469 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1470 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1471 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1472 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1473 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1474 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1475 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd1476 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd1477 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1478 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd1479 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1480 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1481 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1482 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1483 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1484 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1485 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1486 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1487 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd1488 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1489 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd1490 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd1491 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd1492 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd1493 : begin data_real = -16'sd16384; data_imag = 16'sd0; end
		12'd1494 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd1495 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd1496 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd1497 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1498 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd1499 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1500 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1501 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1502 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd1503 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd1504 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1505 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1506 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1507 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1508 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1509 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1510 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1511 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd1512 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1513 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd1514 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1515 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1516 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1517 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1518 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd1519 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd1520 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1521 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1522 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd1523 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1524 : begin data_real = -16'sd14080; data_imag = 16'sd0; end
		12'd1525 : begin data_real = -16'sd18432; data_imag = 16'sd0; end
		12'd1526 : begin data_real = -16'sd16128; data_imag = 16'sd0; end
		12'd1527 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd1528 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd1529 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd1530 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1531 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd1532 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1533 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1534 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd1535 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd1536 : begin data_real = 16'sd18688; data_imag = 16'sd0; end
		12'd1537 : begin data_real = 16'sd16896; data_imag = 16'sd0; end
		12'd1538 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1539 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1540 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1541 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1542 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1543 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1544 : begin data_real = -16'sd16128; data_imag = 16'sd0; end
		12'd1545 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1546 : begin data_real = -16'sd15616; data_imag = 16'sd0; end
		12'd1547 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd1548 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1549 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1550 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1551 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd1552 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd1553 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1554 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1555 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1556 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1557 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1558 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1559 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1560 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1561 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1562 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1563 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd1564 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1565 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1566 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1567 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1568 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd1569 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd1570 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd1571 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd1572 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd1573 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1574 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1575 : begin data_real = -16'sd14336; data_imag = 16'sd0; end
		12'd1576 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1577 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1578 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd1579 : begin data_real = -16'sd22784; data_imag = 16'sd0; end
		12'd1580 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd1581 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd1582 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd1583 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd1584 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1585 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1586 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd1587 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd1588 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd1589 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1590 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd1591 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd1592 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1593 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd1594 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1595 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd1596 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd1597 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1598 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1599 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1600 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1601 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1602 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1603 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1604 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd1605 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd1606 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1607 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd1608 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1609 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1610 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1611 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd1612 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1613 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1614 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1615 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1616 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1617 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1618 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1619 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd1620 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1621 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd1622 : begin data_real = 16'sd13312; data_imag = 16'sd0; end
		12'd1623 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd1624 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd1625 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd1626 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1627 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1628 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1629 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1630 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1631 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd1632 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd1633 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd1634 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1635 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd1636 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1637 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1638 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd1639 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1640 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1641 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd1642 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1643 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1644 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd1645 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1646 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1647 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1648 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1649 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1650 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1651 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1652 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1653 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1654 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1655 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd1656 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd1657 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1658 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1659 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd1660 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1661 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd1662 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1663 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd1664 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1665 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd1666 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd1667 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd1668 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd1669 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd1670 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd1671 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd1672 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd1673 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1674 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1675 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd1676 : begin data_real = 16'sd18944; data_imag = 16'sd0; end
		12'd1677 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1678 : begin data_real = 16'sd16640; data_imag = 16'sd0; end
		12'd1679 : begin data_real = 16'sd16640; data_imag = 16'sd0; end
		12'd1680 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1681 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1682 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd1683 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1684 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1685 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1686 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd1687 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd1688 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1689 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd1690 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd1691 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1692 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1693 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1694 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1695 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1696 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1697 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1698 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1699 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd1700 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1701 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1702 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1703 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd1704 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd1705 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1706 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1707 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1708 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd1709 : begin data_real = 16'sd18688; data_imag = 16'sd0; end
		12'd1710 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1711 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd1712 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd1713 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd1714 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1715 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd1716 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1717 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd1718 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd1719 : begin data_real = -16'sd19456; data_imag = 16'sd0; end
		12'd1720 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd1721 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1722 : begin data_real = -16'sd15872; data_imag = 16'sd0; end
		12'd1723 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd1724 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd1725 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd1726 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd1727 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd1728 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1729 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1730 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd1731 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1732 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd1733 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1734 : begin data_real = 16'sd15104; data_imag = 16'sd0; end
		12'd1735 : begin data_real = 16'sd13312; data_imag = 16'sd0; end
		12'd1736 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1737 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1738 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd1739 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd1740 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1741 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1742 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1743 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd1744 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd1745 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd1746 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1747 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1748 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1749 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1750 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd1751 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd1752 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1753 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd1754 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd1755 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd1756 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1757 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1758 : begin data_real = -16'sd16128; data_imag = 16'sd0; end
		12'd1759 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd1760 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1761 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1762 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd1763 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1764 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd1765 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd1766 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd1767 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1768 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1769 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1770 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1771 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1772 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1773 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1774 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1775 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd1776 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1777 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd1778 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd1779 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1780 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1781 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1782 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1783 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1784 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd1785 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd1786 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd1787 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd1788 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1789 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd1790 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1791 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd1792 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd1793 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1794 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1795 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd1796 : begin data_real = 16'sd15360; data_imag = 16'sd0; end
		12'd1797 : begin data_real = 16'sd17664; data_imag = 16'sd0; end
		12'd1798 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1799 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1800 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd1801 : begin data_real = 16'sd15872; data_imag = 16'sd0; end
		12'd1802 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1803 : begin data_real = 16'sd15360; data_imag = 16'sd0; end
		12'd1804 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd1805 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd1806 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1807 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd1808 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd1809 : begin data_real = -16'sd16128; data_imag = 16'sd0; end
		12'd1810 : begin data_real = -16'sd26112; data_imag = 16'sd0; end
		12'd1811 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1812 : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd1813 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd1814 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1815 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1816 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1817 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd1818 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1819 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1820 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd1821 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd1822 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd1823 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd1824 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1825 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd1826 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1827 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1828 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1829 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1830 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1831 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd1832 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd1833 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1834 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd1835 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1836 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd1837 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1838 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd1839 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1840 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd1841 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd1842 : begin data_real = -16'sd16128; data_imag = 16'sd0; end
		12'd1843 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd1844 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd1845 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1846 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1847 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd1848 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1849 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1850 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd1851 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd1852 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd1853 : begin data_real = 16'sd16896; data_imag = 16'sd0; end
		12'd1854 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd1855 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd1856 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd1857 : begin data_real = 16'sd13312; data_imag = 16'sd0; end
		12'd1858 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1859 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1860 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1861 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd1862 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd1863 : begin data_real = -16'sd16384; data_imag = 16'sd0; end
		12'd1864 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1865 : begin data_real = -16'sd18688; data_imag = 16'sd0; end
		12'd1866 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd1867 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd1868 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd1869 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd1870 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1871 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd1872 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1873 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1874 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1875 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1876 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd1877 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd1878 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd1879 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1880 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1881 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1882 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1883 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd1884 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd1885 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1886 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd1887 : begin data_real = 16'sd17664; data_imag = 16'sd0; end
		12'd1888 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1889 : begin data_real = 16'sd14336; data_imag = 16'sd0; end
		12'd1890 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1891 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd1892 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd1893 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd1894 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd1895 : begin data_real = -16'sd18432; data_imag = 16'sd0; end
		12'd1896 : begin data_real = -16'sd16384; data_imag = 16'sd0; end
		12'd1897 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd1898 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd1899 : begin data_real = -16'sd15616; data_imag = 16'sd0; end
		12'd1900 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1901 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd1902 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd1903 : begin data_real = 16'sd13312; data_imag = 16'sd0; end
		12'd1904 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1905 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1906 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1907 : begin data_real = 16'sd15104; data_imag = 16'sd0; end
		12'd1908 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd1909 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1910 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd1911 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd1912 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1913 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1914 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1915 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd1916 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1917 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1918 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd1919 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd1920 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd1921 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd1922 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd1923 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1924 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1925 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd1926 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1927 : begin data_real = -16'sd17920; data_imag = 16'sd0; end
		12'd1928 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1929 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd1930 : begin data_real = -16'sd17408; data_imag = 16'sd0; end
		12'd1931 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd1932 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1933 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd1934 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1935 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd1936 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd1937 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1938 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd1939 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd1940 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd1941 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd1942 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd1943 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd1944 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd1945 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd1946 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd1947 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd1948 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1949 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1950 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd1951 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd1952 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd1953 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd1954 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd1955 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd1956 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd1957 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd1958 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd1959 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd1960 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd1961 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1962 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd1963 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd1964 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd1965 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd1966 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd1967 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd1968 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd1969 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd1970 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd1971 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd1972 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd1973 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd1974 : begin data_real = 16'sd13312; data_imag = 16'sd0; end
		12'd1975 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd1976 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd1977 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd1978 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1979 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd1980 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd1981 : begin data_real = -16'sd16640; data_imag = 16'sd0; end
		12'd1982 : begin data_real = -16'sd16896; data_imag = 16'sd0; end
		12'd1983 : begin data_real = -16'sd16896; data_imag = 16'sd0; end
		12'd1984 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd1985 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd1986 : begin data_real = -16'sd18688; data_imag = 16'sd0; end
		12'd1987 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd1988 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd1989 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd1990 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd1991 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd1992 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd1993 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd1994 : begin data_real = 16'sd15104; data_imag = 16'sd0; end
		12'd1995 : begin data_real = 16'sd20480; data_imag = 16'sd0; end
		12'd1996 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd1997 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd1998 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd1999 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd2000 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2001 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd2002 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2003 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd2004 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2005 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2006 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2007 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd2008 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2009 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2010 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd2011 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2012 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2013 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2014 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd2015 : begin data_real = -16'sd16896; data_imag = 16'sd0; end
		12'd2016 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2017 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd2018 : begin data_real = -16'sd12032; data_imag = 16'sd0; end
		12'd2019 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2020 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd2021 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd2022 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2023 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2024 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd2025 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2026 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2027 : begin data_real = 16'sd19200; data_imag = 16'sd0; end
		12'd2028 : begin data_real = 16'sd23808; data_imag = 16'sd0; end
		12'd2029 : begin data_real = 16'sd16640; data_imag = 16'sd0; end
		12'd2030 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2031 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd2032 : begin data_real = 16'sd15616; data_imag = 16'sd0; end
		12'd2033 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd2034 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2035 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd2036 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd2037 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd2038 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd2039 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd2040 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2041 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2042 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2043 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2044 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd2045 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2046 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2047 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2048 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2049 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd2050 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2051 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd2052 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2053 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2054 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd2055 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2056 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd2057 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2058 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2059 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2060 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2061 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2062 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd2063 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd2064 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2065 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2066 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2067 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd2068 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd2069 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2070 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd2071 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd2072 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2073 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd2074 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd2075 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd2076 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2077 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd2078 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2079 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2080 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd2081 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd2082 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2083 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2084 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd2085 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2086 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2087 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2088 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd2089 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2090 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd2091 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2092 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd2093 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2094 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2095 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2096 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2097 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2098 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2099 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2100 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2101 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2102 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2103 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2104 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2105 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2106 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2107 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd2108 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd2109 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd2110 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd2111 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd2112 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2113 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2114 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd2115 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd2116 : begin data_real = 16'sd16896; data_imag = 16'sd0; end
		12'd2117 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2118 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2119 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd2120 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2121 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2122 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd2123 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2124 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2125 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2126 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd2127 : begin data_real = -16'sd14080; data_imag = 16'sd0; end
		12'd2128 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2129 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd2130 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2131 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd2132 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2133 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2134 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd2135 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2136 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2137 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd2138 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd2139 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd2140 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2141 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd2142 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2143 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2144 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2145 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd2146 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2147 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2148 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd2149 : begin data_real = 16'sd19200; data_imag = 16'sd0; end
		12'd2150 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2151 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2152 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2153 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd2154 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2155 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2156 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd2157 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd2158 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd2159 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd2160 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2161 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2162 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd2163 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd2164 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd2165 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2166 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd2167 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2168 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2169 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd2170 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2171 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2172 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2173 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd2174 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2175 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2176 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2177 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2178 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd2179 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2180 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd2181 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2182 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2183 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2184 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2185 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2186 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd2187 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2188 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2189 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd2190 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2191 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2192 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd2193 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd2194 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2195 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd2196 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2197 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd2198 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd2199 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2200 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2201 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd2202 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd2203 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd2204 : begin data_real = 16'sd18432; data_imag = 16'sd0; end
		12'd2205 : begin data_real = 16'sd18176; data_imag = 16'sd0; end
		12'd2206 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2207 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2208 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2209 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2210 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2211 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2212 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2213 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2214 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2215 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2216 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2217 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd2218 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd2219 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd2220 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd2221 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd2222 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2223 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd2224 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2225 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2226 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd2227 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd2228 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd2229 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2230 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd2231 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2232 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd2233 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd2234 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2235 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd2236 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd2237 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2238 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd2239 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2240 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2241 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd2242 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2243 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2244 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2245 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2246 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd2247 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd2248 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd2249 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd2250 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd2251 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2252 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd2253 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2254 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd2255 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2256 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2257 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd2258 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd2259 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2260 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2261 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd2262 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2263 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd2264 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2265 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2266 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd2267 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2268 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2269 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2270 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2271 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2272 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2273 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd2274 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd2275 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd2276 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd2277 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2278 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2279 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2280 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd2281 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd2282 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd2283 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd2284 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2285 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd2286 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd2287 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd2288 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd2289 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd2290 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2291 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2292 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2293 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2294 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd2295 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2296 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd2297 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd2298 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2299 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2300 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2301 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2302 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2303 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2304 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd2305 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd2306 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2307 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2308 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd2309 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd2310 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd2311 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2312 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2313 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2314 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2315 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd2316 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd2317 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd2318 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd2319 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd2320 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd2321 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd2322 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd2323 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2324 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2325 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2326 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd2327 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd2328 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd2329 : begin data_real = 16'sd17152; data_imag = 16'sd0; end
		12'd2330 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd2331 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2332 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd2333 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd2334 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2335 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd2336 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2337 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd2338 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd2339 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd2340 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2341 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd2342 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd2343 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2344 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2345 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2346 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2347 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2348 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd2349 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd2350 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2351 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd2352 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2353 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd2354 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd2355 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd2356 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd2357 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2358 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2359 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd2360 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd2361 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd2362 : begin data_real = 16'sd17664; data_imag = 16'sd0; end
		12'd2363 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd2364 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd2365 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2366 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2367 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2368 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd2369 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd2370 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd2371 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd2372 : begin data_real = -16'sd15616; data_imag = 16'sd0; end
		12'd2373 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd2374 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd2375 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd2376 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd2377 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd2378 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2379 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2380 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2381 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd2382 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2383 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd2384 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd2385 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2386 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2387 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2388 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2389 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2390 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd2391 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2392 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2393 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2394 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2395 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd2396 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2397 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2398 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd2399 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd2400 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2401 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2402 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd2403 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2404 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd2405 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd2406 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd2407 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd2408 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2409 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2410 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2411 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2412 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd2413 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2414 : begin data_real = 16'sd24064; data_imag = 16'sd0; end
		12'd2415 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd2416 : begin data_real = 16'sd17152; data_imag = 16'sd0; end
		12'd2417 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2418 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2419 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd2420 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd2421 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2422 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2423 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2424 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd2425 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2426 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2427 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd2428 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd2429 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd2430 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2431 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd2432 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd2433 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2434 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2435 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd2436 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2437 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd2438 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2439 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2440 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2441 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2442 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2443 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2444 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2445 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2446 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd2447 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2448 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd2449 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd2450 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd2451 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd2452 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd2453 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2454 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2455 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd2456 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2457 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd2458 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2459 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd2460 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2461 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd2462 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2463 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2464 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2465 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2466 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd2467 : begin data_real = 16'sd23296; data_imag = 16'sd0; end
		12'd2468 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd2469 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd2470 : begin data_real = 16'sd16384; data_imag = 16'sd0; end
		12'd2471 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd2472 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2473 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd2474 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2475 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd2476 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2477 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2478 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2479 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd2480 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd2481 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd2482 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2483 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd2484 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd2485 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd2486 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd2487 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2488 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd2489 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd2490 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd2491 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2492 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd2493 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd2494 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2495 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd2496 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd2497 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2498 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2499 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2500 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2501 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd2502 : begin data_real = 16'sd18176; data_imag = 16'sd0; end
		12'd2503 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd2504 : begin data_real = 16'sd19200; data_imag = 16'sd0; end
		12'd2505 : begin data_real = 16'sd15104; data_imag = 16'sd0; end
		12'd2506 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd2507 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2508 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2509 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2510 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd2511 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2512 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd2513 : begin data_real = -16'sd18176; data_imag = 16'sd0; end
		12'd2514 : begin data_real = -16'sd16896; data_imag = 16'sd0; end
		12'd2515 : begin data_real = -16'sd14080; data_imag = 16'sd0; end
		12'd2516 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2517 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd2518 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2519 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd2520 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2521 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd2522 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2523 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2524 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2525 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd2526 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2527 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2528 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd2529 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2530 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd2531 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd2532 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2533 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2534 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd2535 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd2536 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2537 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd2538 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd2539 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2540 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd2541 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd2542 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd2543 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd2544 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2545 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd2546 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd2547 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd2548 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd2549 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd2550 : begin data_real = -16'sd15616; data_imag = 16'sd0; end
		12'd2551 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd2552 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd2553 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2554 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd2555 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd2556 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd2557 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd2558 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd2559 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd2560 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd2561 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd2562 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2563 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd2564 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2565 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2566 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd2567 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2568 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd2569 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2570 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2571 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2572 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2573 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2574 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd2575 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2576 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2577 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd2578 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd2579 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2580 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd2581 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd2582 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd2583 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2584 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2585 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2586 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2587 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd2588 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd2589 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd2590 : begin data_real = 16'sd15104; data_imag = 16'sd0; end
		12'd2591 : begin data_real = 16'sd27648; data_imag = 16'sd0; end
		12'd2592 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd2593 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd2594 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2595 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd2596 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd2597 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2598 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2599 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd2600 : begin data_real = -16'sd14336; data_imag = 16'sd0; end
		12'd2601 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd2602 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd2603 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2604 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2605 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2606 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd2607 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2608 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd2609 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2610 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2611 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd2612 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd2613 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd2614 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2615 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd2616 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2617 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2618 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd2619 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2620 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2621 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2622 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2623 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd2624 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd2625 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd2626 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd2627 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd2628 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2629 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2630 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2631 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd2632 : begin data_real = -16'sd14336; data_imag = 16'sd0; end
		12'd2633 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd2634 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2635 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd2636 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd2637 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2638 : begin data_real = -16'sd18176; data_imag = 16'sd0; end
		12'd2639 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd2640 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2641 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2642 : begin data_real = 16'sd17152; data_imag = 16'sd0; end
		12'd2643 : begin data_real = 16'sd14336; data_imag = 16'sd0; end
		12'd2644 : begin data_real = 16'sd17152; data_imag = 16'sd0; end
		12'd2645 : begin data_real = 16'sd15104; data_imag = 16'sd0; end
		12'd2646 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd2647 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd2648 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2649 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2650 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2651 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2652 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2653 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2654 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2655 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd2656 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd2657 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd2658 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2659 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd2660 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2661 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2662 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2663 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2664 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2665 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2666 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2667 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd2668 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd2669 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2670 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd2671 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2672 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2673 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd2674 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2675 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd2676 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd2677 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd2678 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd2679 : begin data_real = 16'sd24320; data_imag = 16'sd0; end
		12'd2680 : begin data_real = 16'sd14336; data_imag = 16'sd0; end
		12'd2681 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2682 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd2683 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2684 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2685 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2686 : begin data_real = -16'sd18176; data_imag = 16'sd0; end
		12'd2687 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2688 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2689 : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd2690 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2691 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd2692 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2693 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd2694 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd2695 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2696 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2697 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2698 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2699 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd2700 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2701 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2702 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2703 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd2704 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd2705 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2706 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd2707 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2708 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2709 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2710 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd2711 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2712 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd2713 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2714 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2715 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2716 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2717 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2718 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2719 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2720 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd2721 : begin data_real = -16'sd18688; data_imag = 16'sd0; end
		12'd2722 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2723 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2724 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd2725 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd2726 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2727 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2728 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2729 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd2730 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd2731 : begin data_real = 16'sd17920; data_imag = 16'sd0; end
		12'd2732 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd2733 : begin data_real = 16'sd16384; data_imag = 16'sd0; end
		12'd2734 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd2735 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2736 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd2737 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd2738 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2739 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd2740 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd2741 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2742 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd2743 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd2744 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd2745 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd2746 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2747 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2748 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2749 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2750 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2751 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2752 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2753 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2754 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2755 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2756 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2757 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2758 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2759 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd2760 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2761 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2762 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd2763 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2764 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd2765 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd2766 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd2767 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd2768 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd2769 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd2770 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2771 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2772 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd2773 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd2774 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd2775 : begin data_real = -16'sd19200; data_imag = 16'sd0; end
		12'd2776 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2777 : begin data_real = -16'sd19456; data_imag = 16'sd0; end
		12'd2778 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd2779 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd2780 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2781 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2782 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2783 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2784 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd2785 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd2786 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd2787 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd2788 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd2789 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd2790 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2791 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd2792 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2793 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd2794 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd2795 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd2796 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2797 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd2798 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd2799 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd2800 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2801 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2802 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2803 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd2804 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd2805 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd2806 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2807 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd2808 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd2809 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd2810 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd2811 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd2812 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd2813 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd2814 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2815 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2816 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2817 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2818 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd2819 : begin data_real = 16'sd15616; data_imag = 16'sd0; end
		12'd2820 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd2821 : begin data_real = 16'sd24064; data_imag = 16'sd0; end
		12'd2822 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2823 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd2824 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd2825 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2826 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2827 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2828 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd2829 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd2830 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd2831 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd2832 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd2833 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd2834 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd2835 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2836 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd2837 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2838 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd2839 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd2840 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2841 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2842 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd2843 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2844 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd2845 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd2846 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2847 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2848 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd2849 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd2850 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2851 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2852 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd2853 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd2854 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd2855 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd2856 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2857 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd2858 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2859 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd2860 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2861 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd2862 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd2863 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2864 : begin data_real = -16'sd14080; data_imag = 16'sd0; end
		12'd2865 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2866 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd2867 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd2868 : begin data_real = -16'sd19200; data_imag = 16'sd0; end
		12'd2869 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd2870 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd2871 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2872 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2873 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd2874 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd2875 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd2876 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd2877 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd2878 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd2879 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd2880 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd2881 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd2882 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd2883 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2884 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd2885 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2886 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2887 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd2888 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2889 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2890 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2891 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2892 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd2893 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd2894 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2895 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd2896 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2897 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd2898 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd2899 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2900 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2901 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd2902 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2903 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd2904 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd2905 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd2906 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2907 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd2908 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd2909 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd2910 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd2911 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd2912 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd2913 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2914 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2915 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2916 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2917 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2918 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd2919 : begin data_real = -16'sd19200; data_imag = 16'sd0; end
		12'd2920 : begin data_real = -16'sd12032; data_imag = 16'sd0; end
		12'd2921 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2922 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2923 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2924 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2925 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd2926 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2927 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd2928 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2929 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd2930 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd2931 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2932 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd2933 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd2934 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2935 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd2936 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd2937 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2938 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2939 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2940 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd2941 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd2942 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd2943 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd2944 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd2945 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2946 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd2947 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2948 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2949 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd2950 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd2951 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd2952 : begin data_real = -16'sd21504; data_imag = 16'sd0; end
		12'd2953 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd2954 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2955 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd2956 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd2957 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd2958 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2959 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd2960 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd2961 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd2962 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd2963 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd2964 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd2965 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd2966 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd2967 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd2968 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd2969 : begin data_real = -16'sd15872; data_imag = 16'sd0; end
		12'd2970 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd2971 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd2972 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd2973 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd2974 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd2975 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd2976 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd2977 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2978 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd2979 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd2980 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd2981 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd2982 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd2983 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd2984 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2985 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd2986 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd2987 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd2988 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd2989 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd2990 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd2991 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd2992 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd2993 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd2994 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd2995 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd2996 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd2997 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd2998 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd2999 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3000 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3001 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3002 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3003 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd3004 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd3005 : begin data_real = -16'sd15872; data_imag = 16'sd0; end
		12'd3006 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd3007 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd3008 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd3009 : begin data_real = -16'sd15616; data_imag = 16'sd0; end
		12'd3010 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3011 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3012 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd3013 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3014 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3015 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd3016 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3017 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3018 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3019 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd3020 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3021 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3022 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3023 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd3024 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3025 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3026 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3027 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3028 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd3029 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3030 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd3031 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd3032 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd3033 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd3034 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3035 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3036 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd3037 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd3038 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3039 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3040 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3041 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3042 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3043 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3044 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd3045 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3046 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3047 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3048 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3049 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd3050 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd3051 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd3052 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3053 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3054 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd3055 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd3056 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3057 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3058 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3059 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3060 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3061 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3062 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3063 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3064 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd3065 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3066 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3067 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd3068 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3069 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3070 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd3071 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3072 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3073 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3074 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3075 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd3076 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd3077 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3078 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3079 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3080 : begin data_real = 16'sd14336; data_imag = 16'sd0; end
		12'd3081 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd3082 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd3083 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3084 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd3085 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3086 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3087 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3088 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd3089 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd3090 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3091 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3092 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3093 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3094 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd3095 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3096 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd3097 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3098 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd3099 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3100 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd3101 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3102 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3103 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3104 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd3105 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3106 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3107 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3108 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3109 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3110 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3111 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd3112 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd3113 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3114 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3115 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd3116 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd3117 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd3118 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd3119 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3120 : begin data_real = 16'sd18688; data_imag = 16'sd0; end
		12'd3121 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3122 : begin data_real = 16'sd15360; data_imag = 16'sd0; end
		12'd3123 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd3124 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3125 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3126 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3127 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd3128 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd3129 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3130 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3131 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3132 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3133 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3134 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3135 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3136 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd3137 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd3138 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd3139 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3140 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3141 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3142 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd3143 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3144 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd3145 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd3146 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3147 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd3148 : begin data_real = -16'sd18176; data_imag = 16'sd0; end
		12'd3149 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3150 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3151 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3152 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd3153 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3154 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd3155 : begin data_real = 16'sd14080; data_imag = 16'sd0; end
		12'd3156 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3157 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3158 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3159 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3160 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3161 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd3162 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3163 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3164 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3165 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3166 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3167 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd3168 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3169 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3170 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd3171 : begin data_real = 16'sd15872; data_imag = 16'sd0; end
		12'd3172 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd3173 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd3174 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd3175 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3176 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd3177 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3178 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd3179 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3180 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3181 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3182 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3183 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3184 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3185 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3186 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3187 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3188 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd3189 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd3190 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3191 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3192 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3193 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3194 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3195 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3196 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd3197 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3198 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3199 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3200 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3201 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3202 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd3203 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd3204 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd3205 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3206 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3207 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd3208 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd3209 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd3210 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3211 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3212 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd3213 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3214 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3215 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3216 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3217 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd3218 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3219 : begin data_real = -16'sd18432; data_imag = 16'sd0; end
		12'd3220 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3221 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3222 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3223 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3224 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3225 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3226 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3227 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3228 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3229 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd3230 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd3231 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3232 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd3233 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3234 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd3235 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3236 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3237 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd3238 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3239 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3240 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3241 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3242 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd3243 : begin data_real = 16'sd22528; data_imag = 16'sd0; end
		12'd3244 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd3245 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3246 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3247 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3248 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3249 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd3250 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd3251 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3252 : begin data_real = -16'sd18944; data_imag = 16'sd0; end
		12'd3253 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3254 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd3255 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd3256 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3257 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3258 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3259 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd3260 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd3261 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3262 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3263 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3264 : begin data_real = 16'sd12032; data_imag = 16'sd0; end
		12'd3265 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3266 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3267 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd3268 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3269 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3270 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd3271 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd3272 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd3273 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3274 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd3275 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3276 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd3277 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd3278 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3279 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3280 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd3281 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd3282 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd3283 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd3284 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd3285 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3286 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd3287 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd3288 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd3289 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3290 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3291 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd3292 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd3293 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3294 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd3295 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd3296 : begin data_real = 16'sd16384; data_imag = 16'sd0; end
		12'd3297 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd3298 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd3299 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3300 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd3301 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd3302 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3303 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3304 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd3305 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3306 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd3307 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3308 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3309 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3310 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd3311 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd3312 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3313 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3314 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd3315 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3316 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3317 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd3318 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3319 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd3320 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd3321 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3322 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3323 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3324 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd3325 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3326 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3327 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3328 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3329 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd3330 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd3331 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3332 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3333 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3334 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd3335 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3336 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd3337 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd3338 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd3339 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3340 : begin data_real = -16'sd18944; data_imag = 16'sd0; end
		12'd3341 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3342 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd3343 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3344 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3345 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3346 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3347 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3348 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd3349 : begin data_real = 16'sd17920; data_imag = 16'sd0; end
		12'd3350 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd3351 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd3352 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3353 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3354 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3355 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3356 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3357 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3358 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3359 : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd3360 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd3361 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3362 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3363 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd3364 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd3365 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3366 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3367 : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd3368 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3369 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd3370 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3371 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd3372 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3373 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd3374 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3375 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3376 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3377 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3378 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3379 : begin data_real = 16'sd14336; data_imag = 16'sd0; end
		12'd3380 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd3381 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd3382 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd3383 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd3384 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd3385 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd3386 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd3387 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd3388 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3389 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3390 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd3391 : begin data_real = -16'sd16640; data_imag = 16'sd0; end
		12'd3392 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd3393 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd3394 : begin data_real = -16'sd19200; data_imag = 16'sd0; end
		12'd3395 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd3396 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3397 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd3398 : begin data_real = -16'sd10752; data_imag = 16'sd0; end
		12'd3399 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3400 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3401 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3402 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3403 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd3404 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd3405 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd3406 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd3407 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3408 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3409 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3410 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3411 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3412 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3413 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd3414 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3415 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd3416 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3417 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd3418 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3419 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3420 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3421 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3422 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3423 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd3424 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3425 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3426 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd3427 : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd3428 : begin data_real = -16'sd18176; data_imag = 16'sd0; end
		12'd3429 : begin data_real = -16'sd12032; data_imag = 16'sd0; end
		12'd3430 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3431 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd3432 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3433 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3434 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd3435 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd3436 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd3437 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd3438 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3439 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd3440 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3441 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3442 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3443 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd3444 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3445 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd3446 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3447 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd3448 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3449 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3450 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3451 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3452 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3453 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3454 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3455 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd3456 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3457 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3458 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd3459 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd3460 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd3461 : begin data_real = -16'sd14080; data_imag = 16'sd0; end
		12'd3462 : begin data_real = -16'sd11008; data_imag = 16'sd0; end
		12'd3463 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3464 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd3465 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3466 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3467 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd3468 : begin data_real = 16'sd13312; data_imag = 16'sd0; end
		12'd3469 : begin data_real = 16'sd18944; data_imag = 16'sd0; end
		12'd3470 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd3471 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd3472 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd3473 : begin data_real = 16'sd19200; data_imag = 16'sd0; end
		12'd3474 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3475 : begin data_real = 16'sd21248; data_imag = 16'sd0; end
		12'd3476 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3477 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3478 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3479 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3480 : begin data_real = -16'sd15872; data_imag = 16'sd0; end
		12'd3481 : begin data_real = -16'sd15616; data_imag = 16'sd0; end
		12'd3482 : begin data_real = -16'sd15616; data_imag = 16'sd0; end
		12'd3483 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3484 : begin data_real = -16'sd16128; data_imag = 16'sd0; end
		12'd3485 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3486 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3487 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3488 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3489 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3490 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd3491 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3492 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd3493 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3494 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3495 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd3496 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3497 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd3498 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd3499 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3500 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3501 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd3502 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3503 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd3504 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3505 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd3506 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3507 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd3508 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3509 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd3510 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3511 : begin data_real = -16'sd16640; data_imag = 16'sd0; end
		12'd3512 : begin data_real = -16'sd14336; data_imag = 16'sd0; end
		12'd3513 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd3514 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd3515 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd3516 : begin data_real = -16'sd11264; data_imag = 16'sd0; end
		12'd3517 : begin data_real = -16'sd9472; data_imag = 16'sd0; end
		12'd3518 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3519 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3520 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3521 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd3522 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3523 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd3524 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd3525 : begin data_real = 16'sd18432; data_imag = 16'sd0; end
		12'd3526 : begin data_real = 16'sd13312; data_imag = 16'sd0; end
		12'd3527 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3528 : begin data_real = 16'sd13824; data_imag = 16'sd0; end
		12'd3529 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd3530 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3531 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd3532 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd3533 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3534 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd3535 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd3536 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd3537 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3538 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3539 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3540 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3541 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3542 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3543 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3544 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd3545 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3546 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3547 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3548 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd3549 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd3550 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd3551 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3552 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3553 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3554 : begin data_real = 16'sd10752; data_imag = 16'sd0; end
		12'd3555 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd3556 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3557 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd3558 : begin data_real = 16'sd11520; data_imag = 16'sd0; end
		12'd3559 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd3560 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3561 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3562 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3563 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3564 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd3565 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3566 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd3567 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd3568 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3569 : begin data_real = -16'sd19200; data_imag = 16'sd0; end
		12'd3570 : begin data_real = -16'sd17920; data_imag = 16'sd0; end
		12'd3571 : begin data_real = -16'sd25856; data_imag = 16'sd0; end
		12'd3572 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3573 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd3574 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3575 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3576 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3577 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd3578 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd3579 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd3580 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3581 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3582 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd3583 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3584 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3585 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3586 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd3587 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3588 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3589 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3590 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3591 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3592 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3593 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3594 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3595 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3596 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3597 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3598 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3599 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3600 : begin data_real = -16'sd17664; data_imag = 16'sd0; end
		12'd3601 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd3602 : begin data_real = -16'sd17152; data_imag = 16'sd0; end
		12'd3603 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd3604 : begin data_real = -16'sd10496; data_imag = 16'sd0; end
		12'd3605 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd3606 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd3607 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd3608 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3609 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd3610 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd3611 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd3612 : begin data_real = 16'sd17152; data_imag = 16'sd0; end
		12'd3613 : begin data_real = 16'sd21248; data_imag = 16'sd0; end
		12'd3614 : begin data_real = 16'sd19968; data_imag = 16'sd0; end
		12'd3615 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3616 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3617 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3618 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd3619 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3620 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd3621 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3622 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3623 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3624 : begin data_real = -16'sd16384; data_imag = 16'sd0; end
		12'd3625 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd3626 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd3627 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3628 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3629 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3630 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3631 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3632 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd3633 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3634 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3635 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3636 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd3637 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd3638 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd3639 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3640 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3641 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd3642 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3643 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3644 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd3645 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd3646 : begin data_real = 16'sd10240; data_imag = 16'sd0; end
		12'd3647 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3648 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3649 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd3650 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3651 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3652 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3653 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd3654 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd3655 : begin data_real = -16'sd18688; data_imag = 16'sd0; end
		12'd3656 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd3657 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd3658 : begin data_real = -16'sd14592; data_imag = 16'sd0; end
		12'd3659 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3660 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3661 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3662 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd3663 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd3664 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd3665 : begin data_real = 16'sd13568; data_imag = 16'sd0; end
		12'd3666 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd3667 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd3668 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd3669 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3670 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3671 : begin data_real = 16'sd12544; data_imag = 16'sd0; end
		12'd3672 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3673 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3674 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd3675 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3676 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3677 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3678 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3679 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3680 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3681 : begin data_real = 16'sd6912; data_imag = 16'sd0; end
		12'd3682 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3683 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd3684 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3685 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3686 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3687 : begin data_real = -16'sd19456; data_imag = 16'sd0; end
		12'd3688 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3689 : begin data_real = -16'sd16896; data_imag = 16'sd0; end
		12'd3690 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd3691 : begin data_real = -16'sd9728; data_imag = 16'sd0; end
		12'd3692 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd3693 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3694 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd3695 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3696 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd3697 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3698 : begin data_real = 16'sd14848; data_imag = 16'sd0; end
		12'd3699 : begin data_real = 16'sd11264; data_imag = 16'sd0; end
		12'd3700 : begin data_real = 16'sd24320; data_imag = 16'sd0; end
		12'd3701 : begin data_real = 16'sd15104; data_imag = 16'sd0; end
		12'd3702 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3703 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd3704 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3705 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3706 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3707 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3708 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3709 : begin data_real = -16'sd20992; data_imag = 16'sd0; end
		12'd3710 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd3711 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd3712 : begin data_real = -16'sd13824; data_imag = 16'sd0; end
		12'd3713 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd3714 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd3715 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3716 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd3717 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3718 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3719 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3720 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3721 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3722 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd3723 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3724 : begin data_real = -16'sd11776; data_imag = 16'sd0; end
		12'd3725 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3726 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3727 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3728 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3729 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3730 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3731 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd3732 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd3733 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3734 : begin data_real = 16'sd17664; data_imag = 16'sd0; end
		12'd3735 : begin data_real = 16'sd16384; data_imag = 16'sd0; end
		12'd3736 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd3737 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3738 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3739 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3740 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd3741 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3742 : begin data_real = -16'sd14080; data_imag = 16'sd0; end
		12'd3743 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3744 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3745 : begin data_real = -16'sd15104; data_imag = 16'sd0; end
		12'd3746 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd3747 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3748 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd3749 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd3750 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3751 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3752 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3753 : begin data_real = 16'sd16384; data_imag = 16'sd0; end
		12'd3754 : begin data_real = 16'sd14336; data_imag = 16'sd0; end
		12'd3755 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3756 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd3757 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3758 : begin data_real = 16'sd2560; data_imag = 16'sd0; end
		12'd3759 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd3760 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3761 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3762 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3763 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3764 : begin data_real = 16'sd5120; data_imag = 16'sd0; end
		12'd3765 : begin data_real = -16'sd2560; data_imag = 16'sd0; end
		12'd3766 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd3767 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3768 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd3769 : begin data_real = 16'sd512; data_imag = 16'sd0; end
		12'd3770 : begin data_real = 16'sd2816; data_imag = 16'sd0; end
		12'd3771 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3772 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3773 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3774 : begin data_real = -16'sd3584; data_imag = 16'sd0; end
		12'd3775 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3776 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3777 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd3778 : begin data_real = -16'sd12032; data_imag = 16'sd0; end
		12'd3779 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3780 : begin data_real = -16'sd8448; data_imag = 16'sd0; end
		12'd3781 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd3782 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd3783 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3784 : begin data_real = 16'sd13312; data_imag = 16'sd0; end
		12'd3785 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3786 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd3787 : begin data_real = 16'sd18176; data_imag = 16'sd0; end
		12'd3788 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd3789 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd3790 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd3791 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3792 : begin data_real = 16'sd17408; data_imag = 16'sd0; end
		12'd3793 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3794 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3795 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3796 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3797 : begin data_real = -16'sd12800; data_imag = 16'sd0; end
		12'd3798 : begin data_real = -16'sd16128; data_imag = 16'sd0; end
		12'd3799 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3800 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd3801 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3802 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3803 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd3804 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3805 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3806 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3807 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd3808 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3809 : begin data_real = 16'sd2048; data_imag = 16'sd0; end
		12'd3810 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3811 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3812 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3813 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3814 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3815 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3816 : begin data_real = -16'sd7680; data_imag = 16'sd0; end
		12'd3817 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd3818 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3819 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3820 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3821 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd3822 : begin data_real = 16'sd11776; data_imag = 16'sd0; end
		12'd3823 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3824 : begin data_real = 16'sd15616; data_imag = 16'sd0; end
		12'd3825 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3826 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3827 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3828 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd3829 : begin data_real = -16'sd7424; data_imag = 16'sd0; end
		12'd3830 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3831 : begin data_real = -16'sd10240; data_imag = 16'sd0; end
		12'd3832 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd3833 : begin data_real = -16'sd19712; data_imag = 16'sd0; end
		12'd3834 : begin data_real = -16'sd8704; data_imag = 16'sd0; end
		12'd3835 : begin data_real = -16'sd11520; data_imag = 16'sd0; end
		12'd3836 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3837 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3838 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3839 : begin data_real = 16'sd1536; data_imag = 16'sd0; end
		12'd3840 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd3841 : begin data_real = 16'sd7936; data_imag = 16'sd0; end
		12'd3842 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3843 : begin data_real = -16'sd3840; data_imag = 16'sd0; end
		12'd3844 : begin data_real = 16'sd4864; data_imag = 16'sd0; end
		12'd3845 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3846 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3847 : begin data_real = 16'sd256; data_imag = 16'sd0; end
		12'd3848 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3849 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3850 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3851 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd3852 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3853 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd3854 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3855 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3856 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3857 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd3858 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3859 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3860 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd3861 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3862 : begin data_real = -16'sd13056; data_imag = 16'sd0; end
		12'd3863 : begin data_real = -16'sd1536; data_imag = 16'sd0; end
		12'd3864 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd3865 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3866 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3867 : begin data_real = -16'sd5120; data_imag = 16'sd0; end
		12'd3868 : begin data_real = -16'sd15360; data_imag = 16'sd0; end
		12'd3869 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3870 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3871 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3872 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3873 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3874 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3875 : begin data_real = 16'sd11008; data_imag = 16'sd0; end
		12'd3876 : begin data_real = 16'sd14592; data_imag = 16'sd0; end
		12'd3877 : begin data_real = 16'sd12288; data_imag = 16'sd0; end
		12'd3878 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3879 : begin data_real = 16'sd13056; data_imag = 16'sd0; end
		12'd3880 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3881 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3882 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd3883 : begin data_real = -16'sd7936; data_imag = 16'sd0; end
		12'd3884 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd3885 : begin data_real = -16'sd14848; data_imag = 16'sd0; end
		12'd3886 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3887 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3888 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3889 : begin data_real = -16'sd3328; data_imag = 16'sd0; end
		12'd3890 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd3891 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd3892 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3893 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd3894 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3895 : begin data_real = 16'sd5376; data_imag = 16'sd0; end
		12'd3896 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3897 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3898 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3899 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3900 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3901 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd3902 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3903 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3904 : begin data_real = -16'sd2816; data_imag = 16'sd0; end
		12'd3905 : begin data_real = -16'sd7168; data_imag = 16'sd0; end
		12'd3906 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3907 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3908 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3909 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd3910 : begin data_real = 16'sd2304; data_imag = 16'sd0; end
		12'd3911 : begin data_real = 16'sd6656; data_imag = 16'sd0; end
		12'd3912 : begin data_real = 16'sd18176; data_imag = 16'sd0; end
		12'd3913 : begin data_real = 16'sd9984; data_imag = 16'sd0; end
		12'd3914 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd3915 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3916 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3917 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3918 : begin data_real = -16'sd8192; data_imag = 16'sd0; end
		12'd3919 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd3920 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3921 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3922 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3923 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd3924 : begin data_real = -16'sd12544; data_imag = 16'sd0; end
		12'd3925 : begin data_real = 16'sd3328; data_imag = 16'sd0; end
		12'd3926 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3927 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3928 : begin data_real = 16'sd9472; data_imag = 16'sd0; end
		12'd3929 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3930 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd3931 : begin data_real = -16'sd3072; data_imag = 16'sd0; end
		12'd3932 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3933 : begin data_real = 16'sd5632; data_imag = 16'sd0; end
		12'd3934 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3935 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3936 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd3937 : begin data_real = -16'sd6400; data_imag = 16'sd0; end
		12'd3938 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd3939 : begin data_real = -16'sd512; data_imag = 16'sd0; end
		12'd3940 : begin data_real = -16'sd4608; data_imag = 16'sd0; end
		12'd3941 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3942 : begin data_real = -16'sd6912; data_imag = 16'sd0; end
		12'd3943 : begin data_real = 16'sd1280; data_imag = 16'sd0; end
		12'd3944 : begin data_real = 16'sd3072; data_imag = 16'sd0; end
		12'd3945 : begin data_real = 16'sd8192; data_imag = 16'sd0; end
		12'd3946 : begin data_real = 16'sd9216; data_imag = 16'sd0; end
		12'd3947 : begin data_real = 16'sd7680; data_imag = 16'sd0; end
		12'd3948 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3949 : begin data_real = 16'sd4608; data_imag = 16'sd0; end
		12'd3950 : begin data_real = 16'sd4096; data_imag = 16'sd0; end
		12'd3951 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3952 : begin data_real = -16'sd9984; data_imag = 16'sd0; end
		12'd3953 : begin data_real = 16'sd768; data_imag = 16'sd0; end
		12'd3954 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3955 : begin data_real = -16'sd9216; data_imag = 16'sd0; end
		12'd3956 : begin data_real = -16'sd13568; data_imag = 16'sd0; end
		12'd3957 : begin data_real = -16'sd1024; data_imag = 16'sd0; end
		12'd3958 : begin data_real = -16'sd13312; data_imag = 16'sd0; end
		12'd3959 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3960 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3961 : begin data_real = 16'sd10496; data_imag = 16'sd0; end
		12'd3962 : begin data_real = 16'sd12800; data_imag = 16'sd0; end
		12'd3963 : begin data_real = 16'sd6400; data_imag = 16'sd0; end
		12'd3964 : begin data_real = 16'sd1792; data_imag = 16'sd0; end
		12'd3965 : begin data_real = 16'sd6144; data_imag = 16'sd0; end
		12'd3966 : begin data_real = 16'sd9728; data_imag = 16'sd0; end
		12'd3967 : begin data_real = 16'sd8704; data_imag = 16'sd0; end
		12'd3968 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd3969 : begin data_real = -16'sd256; data_imag = 16'sd0; end
		12'd3970 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3971 : begin data_real = -16'sd2304; data_imag = 16'sd0; end
		12'd3972 : begin data_real = -16'sd6144; data_imag = 16'sd0; end
		12'd3973 : begin data_real = -16'sd8960; data_imag = 16'sd0; end
		12'd3974 : begin data_real = -16'sd6656; data_imag = 16'sd0; end
		12'd3975 : begin data_real = -16'sd5888; data_imag = 16'sd0; end
		12'd3976 : begin data_real = -16'sd1280; data_imag = 16'sd0; end
		12'd3977 : begin data_real = -16'sd5376; data_imag = 16'sd0; end
		12'd3978 : begin data_real = 16'sd16640; data_imag = 16'sd0; end
		12'd3979 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3980 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3981 : begin data_real = 16'sd3584; data_imag = 16'sd0; end
		12'd3982 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd3983 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3984 : begin data_real = -16'sd5632; data_imag = 16'sd0; end
		12'd3985 : begin data_real = 16'sd4352; data_imag = 16'sd0; end
		12'd3986 : begin data_real = 16'sd5888; data_imag = 16'sd0; end
		12'd3987 : begin data_real = -16'sd4352; data_imag = 16'sd0; end
		12'd3988 : begin data_real = 16'sd1024; data_imag = 16'sd0; end
		12'd3989 : begin data_real = -16'sd4096; data_imag = 16'sd0; end
		12'd3990 : begin data_real = -16'sd12288; data_imag = 16'sd0; end
		12'd3991 : begin data_real = -16'sd768; data_imag = 16'sd0; end
		12'd3992 : begin data_real = -16'sd4864; data_imag = 16'sd0; end
		12'd3993 : begin data_real = -16'sd1792; data_imag = 16'sd0; end
		12'd3994 : begin data_real = -16'sd2048; data_imag = 16'sd0; end
		12'd3995 : begin data_real = 16'sd8448; data_imag = 16'sd0; end
		12'd3996 : begin data_real = 16'sd8960; data_imag = 16'sd0; end
		12'd3997 : begin data_real = 16'sd3840; data_imag = 16'sd0; end
		12'd3998 : begin data_real = 16'sd7168; data_imag = 16'sd0; end
		12'd3999 : begin data_real = 16'sd7424; data_imag = 16'sd0; end
		12'd4000 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4001 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4002 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4003 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4004 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4005 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4006 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4007 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4008 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4009 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4010 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4011 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4012 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4013 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4014 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4015 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4016 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4017 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4018 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4019 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4020 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4021 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4022 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4023 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4024 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4025 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4026 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4027 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4028 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4029 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4030 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4031 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4032 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4033 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4034 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4035 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4036 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4037 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4038 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4039 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4040 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4041 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4042 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4043 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4044 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4045 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4046 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4047 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4048 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4049 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4050 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4051 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4052 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4053 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4054 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4055 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4056 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4057 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4058 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4059 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4060 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4061 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4062 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4063 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4064 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4065 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4066 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4067 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4068 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4069 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4070 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4071 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4072 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4073 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4074 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4075 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4076 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4077 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4078 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4079 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4080 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4081 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4082 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4083 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4084 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4085 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4086 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4087 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4088 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4089 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4090 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4091 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4092 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4093 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4094 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		12'd4095 : begin data_real = 16'sd0; data_imag = 16'sd0; end
		default: begin data_real = 16'sd0; data_imag = 16'sd0; end
        endcase
    end
endmodule

